
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity muxRegFile32x1 is
PORT(	I0: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I1: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I2: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I3: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I4: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I5: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I6: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I7: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I8: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I9: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I10: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I11: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I12: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I13: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I14: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I15: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I16: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I17: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I18: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I19: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I20: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I21: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I22: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I23: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I24: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I25: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I26: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I27: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I28: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I29: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I30: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		I31: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		S:	IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		O:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
end muxRegFile32x1;

architecture Behavioral of muxRegFile32x1 is

begin
O <= 	I0 when  S="00000" else 
		I1 when  S="00001" else 
		I2 when  S="00010" else 
		I3 when  S="00011" else 
		I4 when  S="00100" else 
		I5 when  S="00101" else 
		I6 when  S="00110" else 
		I7 when  S="00111" else 
		I8 when  S="01000" else 
		I9 when  S="01001" else 
		I10 when S="01010" else 
		I11 when S="01011" else 
		I12 when S="01100" else 
		I13 when S="01101" else 
		I14 when S="01110" else 
		I15 when S="01111" else 
		I16 when S="10000" else 
		I17 when S="10001" else 
		I18 when S="10010" else 
		I19 when S="10011" else 
		I20 when S="10100" else 
		I21 when S="10101" else 
		I22 when S="10110" else 
		I23 when S="10111" else 
		I24 when S="11000" else 
		I25 when S="11001" else 
		I26 when S="11010" else 
		I27 when S="11011" else 
		I28 when S="11100" else 
		I29 when S="11101" else 
		I30 when S="11110" else 
		I31 when S="11111" else 
		"ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ";

end Behavioral;

